`timescale 1ns / 1ps
/**
 *
 * Wrapper module that combines processor with its related elements.
 *
 **/

module ProcWrapper (clock, reset);
	input clock, reset;

	wire rwe, mwe, iwe;
	wire[4:0] rd, rs1, rs2, rs3;
	wire[31:0] instAddr, instData, instDataIn, 
		rData, regA, regB, regC,
		memAddr, memDataIn, memDataOut;
	wire [7:0] buttons;


	// ADD YOUR MEMORY FILE HERE
	localparam INSTR_FILE = "";
	
	// Main Processing Unit
	processor CPU(.clock(clock), .reset(reset), 
		/**	   OLD VERSION WITH MEM FILE				
		// ROM
		.address_imem(instAddr), .q_imem(instData),
		**/

		//instRAM
		.address_imem(insAddr), .q_imem(instData),
		.iwren(iwe), .data_imem(instDataIn),

		// Regfile
		.ctrl_writeEnable(rwe),     .ctrl_writeReg(rd),
		.ctrl_readRegA(rs1),     .ctrl_readRegB(rs2), 
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB),
									
		// RAM
		.wren(mwe), .address_dmem(memAddr), 
		.data(memDataIn), .q_dmem(memDataOut),
		
		// Controller
		.controller(buttons)); 
	
	/**     OLD VERSION WITH MEM FILE
	// Instruction Memory (ROM)
	ROM #(.MEMFILE({INSTR_FILE, ".mem"}))
	InstMem(.clk(clock), 
		.addr(instAddr[11:0]), 
		.dataOut(instData));
	**/

	// Instruction Memory (RAM)
	// read from SD card
	RAM InstMem(.clk(clock),
		.wEn(iwe),
		.addr(instAddr[11:0]),
		.dataIn(instDataIn),
		.dataOut(instData));

	// Register File
	regfile RegisterFile(.clock(clock), 
		.ctrl_writeEnable(rwe), .ctrl_reset(reset), 
		.ctrl_writeReg(rd),
		.ctrl_readRegA(rs1), .ctrl_readRegB(rs2), 
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB));
						
	// Processor Memory (RAM)
	RAM ProcMem(.clk(clock), 
		.wEn(mwe), 
		.addr(memAddr[11:0]), 
		.dataIn(memDataIn), 
		.dataOut(memDataOut));
	
	// for testing purposes, assign the buttons to a constant
	assign buttons = 8'b00100110; // B, Left, and Down

endmodule
