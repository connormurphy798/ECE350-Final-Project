/**
 *
 *  The GuyBox.
 *
 **/

module GuyBox(

    );